// Test class instantiates the environment and starts it.

// 测试实例
class test;

  env e0;  // 环境

  function new();
    e0 = new;
  endfunction

  task run();
    e0.run();
  endtask
endclass
