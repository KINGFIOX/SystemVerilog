// 类型的强制转换

module tb;

  byte unsigned ubyte;
  int si = signed'(ubyte);

endmodule
